module Mux8_4b(S2, S1, S0, W0, W1, W2, W3, W4, W5, W6, W7, F);
 input S2, S1, S0;
 input [3:0] W0, W1, W2, W3, W4, W5, W6, W7;
 output [3:0] F;
 
 assign F[0] = (S2&S1&S0&W7[0]) | (S2&S1&~S0&W6[0]) | (S2&~S1&S0&W5[0]) | (S2&~S1&~S0&W4[0]) | (~S2&S1&S0&W3[0]) | (~S2&S1&~S0&W2[0]) | 
				(~S2&~S1&S0&W1[0]) | (~S2&~S1&~S0&W0[0]);
				
 assign F[1] = (S2&S1&S0&W7[1]) | (S2&S1&~S0&W6[1]) | (S2&~S1&S0&W5[1]) | (S2&~S1&~S0&W4[1]) | (~S2&S1&S0&W3[1]) | (~S2&S1&~S0&W2[1]) | 
				(~S2&~S1&S0&W1[1]) | (~S2&~S1&~S0&W0[1]);
				
 assign F[2] = (S2&S1&S0&W7[2]) | (S2&S1&~S0&W6[2]) | (S2&~S1&S0&W5[2]) | (S2&~S1&~S0&W4[2]) | (~S2&S1&S0&W3[2]) | (~S2&S1&~S0&W2[2]) | 
				(~S2&~S1&S0&W1[2]) | (~S2&~S1&~S0&W0[2]);
				
 assign F[3] = (S2&S1&S0&W7[3]) | (S2&S1&~S0&W6[3]) | (S2&~S1&S0&W5[3]) | (S2&~S1&~S0&W4[3]) | (~S2&S1&S0&W3[3]) | (~S2&S1&~S0&W2[3]) | 
				(~S2&~S1&S0&W1[3]) | (~S2&~S1&~S0&W0[3]);
				

				
endmodule